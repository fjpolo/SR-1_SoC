module ROM16_FP2I (
        output logic [15:0] dout, //output [15:0] dout
        input logic [3:0] ad //input [3:0] ad
    );
	
	logic [15:0] prog_to_load [16] = '{
		'{16'b0000000000000000}, 	//00 A	---------
		'{16'b0000000000000001},	//01 B	|A B C D|
		'{16'b0000000000000010},	//02 C	|E F G H|
		'{16'b0000000000000100},	//03 D	|I J K L|
		'{16'b0000000000001000}, 	//04 E	|M N O P|
		'{16'b0000000000010000}, 	//05 F	---------
		'{16'b0000000000100000},	//06 G
		'{16'b0000000001000000}, 	//07 H
		'{16'b0000000010000000}, 	//08 I
		'{16'b0000000100000000},	//09 J
		'{16'b0000001000000000}, 	//10 K
		'{16'b0000010000000000},	//11 L
		'{16'b0000100000000000}, 	//12 M
		'{16'b0001000000000000}, 	//13 N
		'{16'b0010000000000000}, 	//14 O
		'{16'b0100000000000000} 	//15 P
	};
	
	assign dout = prog_to_load[ad];
	
endmodule