module MULT18 (output logic [35:0] dout, input logic [17:0] a, b);
	assign dout = a * b;
endmodule