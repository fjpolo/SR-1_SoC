package MicrocodePackage;
	typedef enum logic [5:0] {
		ENDMICRO,
		RAM_to_A,
		A_to_B,
		A_to_C,
		A_to_D,
		RAM_to_D,
		RAM_to_IR,
		A_to_RAM,
		B_to_A,
		C_to_A,
		RAM_to_PC,
		RAM_to_PC_CF,
		RAM_to_PC_ZF,
		PC_to_RAM,
		PC_to_MAR,
		PC_to_MAR_ADDR,
		RAM_to_MAR,
		RAM_to_MTAR,
		START_BCD,
		ALU_ADD,
		ALU_SUB,
		ALU_MULT,
		ALU_AND,
		ALU_OR,
		ALU_XOR,
		ALU_NOT,
		ALU_AND_B,
		ALU_OR_B,
		ALU_XOR_B,
		ALU_NOT_B,
		ALU_LSHIFT,
		ALU_RSHIFT,
		HLT_CLK,
		INC_PC,
		SET_HALF,
		SET_FULL,
		WAIT_CYCLE,
		DATA_XFER,
		SET_MTAR_GPU,
		START_MT,
		START_UT,
		WAIT_MT,
		WAIT_UT,
		WAIT_FT,
		WAIT_DD,
		WAIT_GPU,
		START_GPU
	} Microcode_enum;
endpackage