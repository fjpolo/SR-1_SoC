//Copyright (C)2014-2024 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.10.03 Education (64-bit)
//Part Number: GW1NR-LV9QN88PC6/I5
//Device: GW1NR-9
//Device Version: C
//Created Time: Mon Feb 24 16:19:21 2025

module DP_BSRAM (douta, doutb, clka, ocea, cea, reseta, wrea, clkb, oceb, ceb, resetb, wreb, ada, dina, adb, dinb);

output [7:0] douta;
output [7:0] doutb;
input clka;
input ocea;
input cea;
input reseta;
input wrea;
input clkb;
input oceb;
input ceb;
input resetb;
input wreb;
input [10:0] ada;
input [7:0] dina;
input [10:0] adb;
input [7:0] dinb;

wire [7:0] dpb_inst_0_douta_w;
wire [7:0] dpb_inst_0_doutb_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

DPB dpb_inst_0 (
    .DOA({dpb_inst_0_douta_w[7:0],douta[7:0]}),
    .DOB({dpb_inst_0_doutb_w[7:0],doutb[7:0]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,gw_gnd}),
    .BLKSELB({gw_gnd,gw_gnd,gw_gnd}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[7:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[7:0]})
);

defparam dpb_inst_0.READ_MODE0 = 1'b0;
defparam dpb_inst_0.READ_MODE1 = 1'b0;
defparam dpb_inst_0.WRITE_MODE0 = 2'b00;
defparam dpb_inst_0.WRITE_MODE1 = 2'b00;
defparam dpb_inst_0.BIT_WIDTH_0 = 8;
defparam dpb_inst_0.BIT_WIDTH_1 = 8;
defparam dpb_inst_0.BLK_SEL_0 = 3'b000;
defparam dpb_inst_0.BLK_SEL_1 = 3'b000;
defparam dpb_inst_0.RESET_MODE = "ASYNC";
defparam dpb_inst_0.INIT_RAM_00 = 256'h0019800000000000000900000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_01 = 256'h0039900600000000003990000000000000399000000000000039800000000000;
defparam dpb_inst_0.INIT_RAM_02 = 256'h00399F09FC00000000399C0FF80000000039900FE00000000039900F80000000;
defparam dpb_inst_0.INIT_RAM_03 = 256'h003980F804000000003983F80400000000398FF81C00000000399FC87C000000;
defparam dpb_inst_0.INIT_RAM_04 = 256'h00398FFC0000000000399FE00400000000399F800400000000399C3004000000;
defparam dpb_inst_0.INIT_RAM_05 = 256'h003980FBFC0000000039803FF8000000003980FFE0000000003983FF80000000;
defparam dpb_inst_0.INIT_RAM_06 = 256'h003980080400000000399C080400000000399F081C000000003983C8FC000000;
defparam dpb_inst_0.INIT_RAM_07 = 256'h00399FFC1800000000399FE06400000000399F818400000000398C0604000000;
defparam dpb_inst_0.INIT_RAM_08 = 256'h0039900BFC0000000039901FF8000000003990FFE0000000003993FF80000000;
defparam dpb_inst_0.INIT_RAM_09 = 256'h003980C804000000003983080400000000398C081C00000000399008FC000000;
defparam dpb_inst_0.INIT_RAM_0A = 256'h0039800018000000003980006400000000398001840000000039803604000000;
defparam dpb_inst_0.INIT_RAM_0B = 256'h0039800000000000003980000000000000398000000000000039800000000000;
defparam dpb_inst_0.INIT_RAM_0C = 256'h003980007FC00000003980007E00000000398000180000000039800000000000;
defparam dpb_inst_0.INIT_RAM_0D = 256'h0039800061FFE0000039800067FF8000003980007FFE0000003980007FF00000;
defparam dpb_inst_0.INIT_RAM_0E = 256'h0038FFC0600078000039FF006001F8000039F800600FF8000039E000603FF800;
defparam dpb_inst_0.INIT_RAM_0F = 256'h003800FFE0001800003807FFE000180000381FFE6000180000387FF860001800;
defparam dpb_inst_0.INIT_RAM_10 = 256'h0039E00000001800003800018000180000380007E00018000038003FE0001800;
defparam dpb_inst_0.INIT_RAM_11 = 256'h00387FFC000018000039FFE0000018000039FF00000018000039FC0000001800;
defparam dpb_inst_0.INIT_RAM_12 = 256'h0038001FFF800000003800FFFC000000003803FFE000000000381FFF80000000;
defparam dpb_inst_0.INIT_RAM_13 = 256'h003800FFE3FFE0000038003FFFFF800000380007FFFC000000380003FFF00000;
defparam dpb_inst_0.INIT_RAM_14 = 256'h0039FF006000780000387FC06003F80000381FF8600FF800003803FE607FF800;
defparam dpb_inst_0.INIT_RAM_15 = 256'h003800006000180000398000600018000039E000600018000039FC0060001800;
defparam dpb_inst_0.INIT_RAM_16 = 256'h0038000006001800003800001800180000380000600018000038000060001800;
defparam dpb_inst_0.INIT_RAM_17 = 256'h003800008001980000380000000E180000380000003018000038000001C01800;
defparam dpb_inst_0.INIT_RAM_18 = 256'h00380000F000000000380000F000000000380000F000000000380000E0006000;
defparam dpb_inst_0.INIT_RAM_19 = 256'h00380000F000000000380000F000000000380000F000000000380000F0000000;
defparam dpb_inst_0.INIT_RAM_1A = 256'h0039E00010000000003800007000000000380000F000000000380000F0000000;
defparam dpb_inst_0.INIT_RAM_1B = 256'h00387FFC000000000039FFE0000000000039FF00000000000039FC0000000000;
defparam dpb_inst_0.INIT_RAM_1C = 256'h0038801FFF800000003800FFFC000000003803FFE000000000381FFF80000000;
defparam dpb_inst_0.INIT_RAM_1D = 256'h003E000003FFE000003F00001FFF8000003B80007FFC000000398003FFF00000;
defparam dpb_inst_0.INIT_RAM_1E = 256'h0020000000007800003000000003F80000380000000FF800003C0000007FF800;
defparam dpb_inst_0.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

endmodule //DP_BSRAM
