package GPU_MicrocodePackage;
	typedef enum logic [5:0] {
		ENDMICRO_GPU,
		VRAM_to_MAU,
		VRAM_to_MAU_ADD,
		VRAM_to_MRAM,
		MAU_to_VRAM2,
		MAU_to_VRAM4,
		INC_PC_A,
		INC_PC_AB,
		PC_A_to_VMAR_A,
		PC_A_to_VMAR_AB,
		PC_B_to_VMAR_AB,
		PC_AB_to_VMAR_AB,
		CPU_to_VRAM,
		CPU_FP_to_VRAM,
		SEND_FRAME,
		INIT_DISPLAY,
		WAIT_ALL_MAU,
		WAIT_ANY_MAU,
		WAIT_FB,
		WAIT_LDU,
		WAIT_START,
		WAIT_DTCU,
		REPEAT_UCODE,
		CONTINUE_OR_END,
		SET_COLOUR,
		VRAM_to_CPU,
		VRAM_to_FP2I,
		START_MAU4,
		START_MAU2,
		CPU_to_MAT_AD4,
		CPU_to_MAT_AD2,
		PC_A_to_MAT_AD4,
		LOAD_LDU_P0,
		START_LDU,
		DRAW_PIXEL,
		WAIT_CYCLE_GPU,
		CPY_A_to_B
	} GPU_Microcode_enum;
endpackage